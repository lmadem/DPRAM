typedef uvm_sequencer #(packet) sequencer;
