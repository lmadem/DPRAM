//This testplan is to verify the functionality of memory model

//mem_test : The purpose of this test is to verify the basic functionality of the memory design. This includes write operation followed by read operation

//in_order_test : This test includes writing all the address locations in the memory randomly, followed by read operations. This test uses in_order_sequence.sv, custom_scoreboard.sv

//out_of_order_test : This purpose of this test is to perform out of ordering sequence in regards to the address location in the memory. This test uses out_of_order_sequence.sv, out_of_order_scoreboard.sv
